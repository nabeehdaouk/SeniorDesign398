module ff_sync(
	input clk,
	input rst
);
	
endmodule
