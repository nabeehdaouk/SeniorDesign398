module arbiter_tb2();
    

	
	initial begin
	   instr
	end
	
endmodule 
