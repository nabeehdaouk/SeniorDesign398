module top_level_tb;
    
endmodule