module binary_to_gray(
	input clk,
	input rst
);
	
endmodule 
