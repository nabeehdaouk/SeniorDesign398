module async_fifo_top_level(
	input clk,
	input rst
);
	
endmodule
