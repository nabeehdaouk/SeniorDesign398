module gray_to_binary(
	input clk,
	input rst
);
	
endmodule
