module arbiter(
	input clk,
	input rst
);
	
endmodule : arbiter
