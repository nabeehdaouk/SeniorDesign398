module top_level(
    input clk,          //Clock driving design
    input resetn        //Global reset
);
    
endmodule